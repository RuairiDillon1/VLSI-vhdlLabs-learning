LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity t_heartbeat_gen is 
end entity; 

architecture tbench of t_heartbeat_gen is 
begin 

end architecture; 
